// Problem statement
// Build a circuit with no inputs and one output that outputs a constant 0

// Solution: 

module top_module(
	output zero
);
assign zero = 0;
endmodule
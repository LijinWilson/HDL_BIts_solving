// Problem statement
// create a wire (in green) by adding an assign statement to connect in to out

// Solution: 
module top_module( input in, output out );
	assign out = in;
endmodule
// Create a module that implements a NOT gate.

// Solution
module top_module( input in, output out );
	assign out = ~in;
endmodule
